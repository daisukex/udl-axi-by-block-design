// ---------------------------------------------------------------------------
// udl_axi: User design logic
// Copyright 2024 Space Cubics, LLC
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// ---------------------------------------------------------------------------

module udl_axi # (
  parameter CM3SS_UDL_ISR_NUM = 16,
  parameter MAINAXI_UDL_M_AXI_ID_WIDTH = 2,
  parameter MAINAXI_S_AXI_ID_WIDTH = 3
) (
  // System Interface
  input  MAXI_CLK,
  input  REF_CLK,
  input  USER_CLK1,
  input  USER_CLK2,
  input  SYS_RSTB,
  input  SYS_RSTB_SYNC_REFCLK,
  input  SYS_RSTB_SYNC_USERCLK1,
  input  SYS_RSTB_SYNC_USERCLK2,
  input  POR_RSTB,
  input  POR_RSTB_SYNC_REFCLK,
  input  BUS_RSTB,

  output [CM3SS_UDL_ISR_NUM-1:0] UDL_INTISR,

  // UDL AXI4 Master Interface
  output [MAINAXI_UDL_M_AXI_ID_WIDTH-1:0] UDL_AXIM_AWID,
  output [31:0] UDL_AXIM_AWADDR,
  output [7:0] UDL_AXIM_AWLEN,
  output [2:0] UDL_AXIM_AWSIZE,
  output [1:0] UDL_AXIM_AWBURST,
  output UDL_AXIM_AWLOCK,
  output [3:0] UDL_AXIM_AWCACHE,
  output [2:0] UDL_AXIM_AWPROT,
  output [3:0] UDL_AXIM_AWQOS,
  output UDL_AXIM_AWVALID,
  input  UDL_AXIM_AWREADY,
  output [31:0] UDL_AXIM_WDATA,
  output [3:0] UDL_AXIM_WSTRB,
  output UDL_AXIM_WLAST,
  output UDL_AXIM_WVALID,
  input  UDL_AXIM_WREADY,
  input  [MAINAXI_UDL_M_AXI_ID_WIDTH-1:0] UDL_AXIM_BID,
  input  [1:0] UDL_AXIM_BRESP,
  input  UDL_AXIM_BVALID,
  output UDL_AXIM_BREADY,
  output [MAINAXI_UDL_M_AXI_ID_WIDTH-1:0] UDL_AXIM_ARID,
  output [31:0] UDL_AXIM_ARADDR,
  output [7:0] UDL_AXIM_ARLEN,
  output [2:0] UDL_AXIM_ARSIZE,
  output [1:0] UDL_AXIM_ARBURST,
  output UDL_AXIM_ARLOCK,
  output [3:0] UDL_AXIM_ARCACHE,
  output [2:0] UDL_AXIM_ARPROT,
  output [3:0] UDL_AXIM_ARQOS,
  output UDL_AXIM_ARVALID,
  input  UDL_AXIM_ARREADY,
  input  [MAINAXI_UDL_M_AXI_ID_WIDTH-1:0] UDL_AXIM_RID,
  input  [31:0] UDL_AXIM_RDATA,
  input  [1:0] UDL_AXIM_RRESP,
  input  UDL_AXIM_RLAST,
  input  UDL_AXIM_RVALID,
  output UDL_AXIM_RREADY,

  // UDL AXI4 Slave Interface
  input  [MAINAXI_S_AXI_ID_WIDTH-1:0] UDL_AXIS_AWID,
  input  [31:0] UDL_AXIS_AWADDR,
  input  [7:0] UDL_AXIS_AWLEN,
  input  [2:0] UDL_AXIS_AWSIZE,
  input  [1:0] UDL_AXIS_AWBURST,
  input  UDL_AXIS_AWLOCK,
  input  [3:0] UDL_AXIS_AWCACHE,
  input  [2:0] UDL_AXIS_AWPROT,
  input  [3:0] UDL_AXIS_AWREGION,
  input  [3:0] UDL_AXIS_AWQOS,
  input  UDL_AXIS_AWVALID,
  output UDL_AXIS_AWREADY,
  input  [31:0] UDL_AXIS_WDATA,
  input  [3:0] UDL_AXIS_WSTRB,
  input  UDL_AXIS_WLAST,
  input  UDL_AXIS_WVALID,
  output UDL_AXIS_WREADY,
  output [MAINAXI_S_AXI_ID_WIDTH-1:0] UDL_AXIS_BID,
  output [1:0] UDL_AXIS_BRESP,
  output UDL_AXIS_BVALID,
  input  UDL_AXIS_BREADY,
  input  [MAINAXI_S_AXI_ID_WIDTH-1:0] UDL_AXIS_ARID,
  input  [31:0] UDL_AXIS_ARADDR,
  input  [7:0] UDL_AXIS_ARLEN,
  input  [2:0] UDL_AXIS_ARSIZE,
  input  [1:0] UDL_AXIS_ARBURST,
  input  UDL_AXIS_ARLOCK,
  input  [3:0] UDL_AXIS_ARCACHE,
  input  [2:0] UDL_AXIS_ARPROT,
  input  [3:0] UDL_AXIS_ARREGION,
  input  [3:0] UDL_AXIS_ARQOS,
  input  UDL_AXIS_ARVALID,
  output UDL_AXIS_ARREADY,
  output [MAINAXI_S_AXI_ID_WIDTH-1:0] UDL_AXIS_RID,
  output [31:0] UDL_AXIS_RDATA,
  output [1:0] UDL_AXIS_RRESP,
  output UDL_AXIS_RLAST,
  output UDL_AXIS_RVALID,
  input  UDL_AXIS_RREADY,

  // Cortex-M3 JTAG Signals
  output IO_NTRST_I,
  output IO_TDI_I,
  output IO_SWCLKTCK_I,
  output IO_SWDIOTMS_I,
  input  IO_SWDIOTMS_O,
  input  IO_SWDIOTMS_EN,
  input  IO_TDOSWO_O,
  input  IO_TDOSWO_EN,
  input  CM3_UART_TX,
  output CM3_UART_RX,

  // User IO Interface
  (* dont_touch = "yes" *) inout [15:0] UIO1,
  (* dont_touch = "yes" *) inout [15:0] UIO2,
  (* dont_touch = "yes" *) inout [5:0]  UIO4,

  // These signals are mutually connected to the FPGA and TRCH.
  // Their connection paths are determined when ordering the OBC,
  // and it will be implemented in the factory.
  inout [2:0] UIO3,
  inout TRCH_UART_TX,
  inout TRCH_UART_RX,
  inout WDOG_OUT
);

udl_axi_bd udl_axi_bd (
  .MAXI_CLK(MAXI_CLK),
  .REF_CLK(REF_CLK),
  .USER_CLK1(USER_CLK1),
  .USER_CLK2(USER_CLK2),
  .SYS_RSTB(SYS_RSTB),
  .SYS_RSTB_SYNC_REFCLK(SYS_RSTB_SYNC_REFCLK),
  .SYS_RSTB_SYNC_USERCLK1(SYS_RSTB_SYNC_USERCLK1),
  .SYS_RSTB_SYNC_USERCLK2(SYS_RSTB_SYNC_USERCLK2),
  .POR_RSTB(POR_RSTB),
  .POR_RSTB_SYNC_REFCLK(POR_RSTB_SYNC_REFCLK),
  .BUS_RSTB(BUS_RSTB),
  .UDL_INTISR(UDL_INTISR),
  .UDL_AXIM_AWID(UDL_AXIM_AWID),
  .UDL_AXIM_AWADDR(UDL_AXIM_AWADDR),
  .UDL_AXIM_AWLEN(UDL_AXIM_AWLEN),
  .UDL_AXIM_AWSIZE(UDL_AXIM_AWSIZE),
  .UDL_AXIM_AWBURST(UDL_AXIM_AWBURST),
  .UDL_AXIM_AWLOCK(UDL_AXIM_AWLOCK),
  .UDL_AXIM_AWCACHE(UDL_AXIM_AWCACHE),
  .UDL_AXIM_AWPROT(UDL_AXIM_AWPROT),
  .UDL_AXIM_AWQOS(UDL_AXIM_AWQOS),
  .UDL_AXIM_AWVALID(UDL_AXIM_AWVALID),
  .UDL_AXIM_AWREADY(UDL_AXIM_AWREADY),
  .UDL_AXIM_WDATA(UDL_AXIM_WDATA),
  .UDL_AXIM_WSTRB(UDL_AXIM_WSTRB),
  .UDL_AXIM_WLAST(UDL_AXIM_WLAST),
  .UDL_AXIM_WVALID(UDL_AXIM_WVALID),
  .UDL_AXIM_WREADY(UDL_AXIM_WREADY),
  .UDL_AXIM_BID(UDL_AXIM_BID),
  .UDL_AXIM_BRESP(UDL_AXIM_BRESP),
  .UDL_AXIM_BVALID(UDL_AXIM_BVALID),
  .UDL_AXIM_BREADY(UDL_AXIM_BREADY),
  .UDL_AXIM_ARID(UDL_AXIM_ARID),
  .UDL_AXIM_ARADDR(UDL_AXIM_ARADDR),
  .UDL_AXIM_ARLEN(UDL_AXIM_ARLEN),
  .UDL_AXIM_ARSIZE(UDL_AXIM_ARSIZE),
  .UDL_AXIM_ARBURST(UDL_AXIM_ARBURST),
  .UDL_AXIM_ARLOCK(UDL_AXIM_ARLOCK),
  .UDL_AXIM_ARCACHE(UDL_AXIM_ARCACHE),
  .UDL_AXIM_ARPROT(UDL_AXIM_ARPROT),
  .UDL_AXIM_ARQOS(UDL_AXIM_ARQOS),
  .UDL_AXIM_ARVALID(UDL_AXIM_ARVALID),
  .UDL_AXIM_ARREADY(UDL_AXIM_ARREADY),
  .UDL_AXIM_RID(UDL_AXIM_RID),
  .UDL_AXIM_RDATA(UDL_AXIM_RDATA),
  .UDL_AXIM_RRESP(UDL_AXIM_RRESP),
  .UDL_AXIM_RLAST(UDL_AXIM_RLAST),
  .UDL_AXIM_RVALID(UDL_AXIM_RVALID),
  .UDL_AXIM_RREADY(UDL_AXIM_RREADY),
  .UDL_AXIS_AWID(UDL_AXIS_AWID),
  .UDL_AXIS_AWADDR(UDL_AXIS_AWADDR),
  .UDL_AXIS_AWLEN(UDL_AXIS_AWLEN),
  .UDL_AXIS_AWSIZE(UDL_AXIS_AWSIZE),
  .UDL_AXIS_AWBURST(UDL_AXIS_AWBURST),
  .UDL_AXIS_AWLOCK(UDL_AXIS_AWLOCK),
  .UDL_AXIS_AWCACHE(UDL_AXIS_AWCACHE),
  .UDL_AXIS_AWPROT(UDL_AXIS_AWPROT),
  .UDL_AXIS_AWREGION(UDL_AXIS_AWREGION),
  .UDL_AXIS_AWQOS(UDL_AXIS_AWQOS),
  .UDL_AXIS_AWVALID(UDL_AXIS_AWVALID),
  .UDL_AXIS_AWREADY(UDL_AXIS_AWREADY),
  .UDL_AXIS_WDATA(UDL_AXIS_WDATA),
  .UDL_AXIS_WSTRB(UDL_AXIS_WSTRB),
  .UDL_AXIS_WLAST(UDL_AXIS_WLAST),
  .UDL_AXIS_WVALID(UDL_AXIS_WVALID),
  .UDL_AXIS_WREADY(UDL_AXIS_WREADY),
  .UDL_AXIS_BID(UDL_AXIS_BID),
  .UDL_AXIS_BRESP(UDL_AXIS_BRESP),
  .UDL_AXIS_BVALID(UDL_AXIS_BVALID),
  .UDL_AXIS_BREADY(UDL_AXIS_BREADY),
  .UDL_AXIS_ARID(UDL_AXIS_ARID),
  .UDL_AXIS_ARADDR(UDL_AXIS_ARADDR),
  .UDL_AXIS_ARLEN(UDL_AXIS_ARLEN),
  .UDL_AXIS_ARSIZE(UDL_AXIS_ARSIZE),
  .UDL_AXIS_ARBURST(UDL_AXIS_ARBURST),
  .UDL_AXIS_ARLOCK(UDL_AXIS_ARLOCK),
  .UDL_AXIS_ARCACHE(UDL_AXIS_ARCACHE),
  .UDL_AXIS_ARPROT(UDL_AXIS_ARPROT),
  .UDL_AXIS_ARREGION(UDL_AXIS_ARREGION),
  .UDL_AXIS_ARQOS(UDL_AXIS_ARQOS),
  .UDL_AXIS_ARVALID(UDL_AXIS_ARVALID),
  .UDL_AXIS_ARREADY(UDL_AXIS_ARREADY),
  .UDL_AXIS_RID(UDL_AXIS_RID),
  .UDL_AXIS_RDATA(UDL_AXIS_RDATA),
  .UDL_AXIS_RRESP(UDL_AXIS_RRESP),
  .UDL_AXIS_RLAST(UDL_AXIS_RLAST),
  .UDL_AXIS_RVALID(UDL_AXIS_RVALID),
  .UDL_AXIS_RREADY(UDL_AXIS_RREADY),
  .IO_NTRST_I(IO_NTRST_I),
  .IO_TDI_I(IO_TDI_I),
  .IO_SWCLKTCK_I(IO_SWCLKTCK_I),
  .IO_SWDIOTMS_I(IO_SWDIOTMS_I),
  .IO_SWDIOTMS_O(IO_SWDIOTMS_O),
  .IO_SWDIOTMS_EN(IO_SWDIOTMS_EN),
  .IO_TDOSWO_O(IO_TDOSWO_O),
  .IO_TDOSWO_EN(IO_TDOSWO_EN),
  .CM3_UART_TX(CM3_UART_TX),
  .CM3_UART_RX(CM3_UART_RX),
  .UIO1(UIO1),
  .UIO2(UIO2),
  .UIO4(UIO4),
  .UIO3(UIO3),
  .TRCH_UART_TX(TRCH_UART_TX),
  .TRCH_UART_RX(TRCH_UART_RX),
  .WDOG_OUT(WDOG_OUT)
);

endmodule
